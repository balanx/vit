module test2 (

input  [3:0] a1, a2, a3,
input        b1, b2, b3,
input  [7:0] d,
input        e,

output  [263:10] f1, f2, f3160,
output           g1, g2, g3,
output  [7:0] h,
output        j

);

reg [3:0] tmp;

main code will be ignore !

endmodule
