
module  test8 ();


endmodule

module  test9;

parameter   DEVICE_ID  = 16'h0466;
parameter   REV        = 16'hF410;

endmodule
